`timescale 1 ns / 100 ps
`define TESTVECS 8

module tb_array
    reg clk, reset;
    reg [2:0] din, dout;
    
